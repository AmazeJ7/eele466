library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity newtons is
    port(newtons_input : in  std_logic_vector (35 downto 0);
         y 	       : out std_logic_vector (35 downto 0));
end entity;

architecture rsr_arch of rsr is

  begin

end architecture;
